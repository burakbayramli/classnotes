
.TITLE Ornek #1

Vin 0 1 AC 1
R1  1 2 1K
R2  0 2 1K
C1  0 2 1UF

.OPTION OUT=80
.PRINT OP Iter(0) V(2)

.PLOT AC  VDB(2)(-20,0)

.AC 5 1K OCT
